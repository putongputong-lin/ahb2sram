../dv/sramc_if.sv
../dv/sramc_dv_class.sv
../dv/tb_top.sv

../de/ahb2sram.v
../de/sram.v
../de/sram_core.v
../de/sramc_slave.v
